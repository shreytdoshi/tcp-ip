��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�M�N��.��	F(�
��_i�5�O2H��Lj�����;�%�X�aK���0R��E瑊�2�k�P�����*�!d�������YV�LE��Â8��hXl��A Y[��N.	���V1[ �/����*+^�xJ�M�D����r|��V�uF�}x_B���hn�|RK����*����`����V��7�}}�=�B��Z�ٻI�+�k%'�Y$�^��H/`C=��}>r���|���֦�^o���(�M�N��v*c�g��\5F�9�Y��{���k���6���5�.*~d��;�2[�^f�;�y��FXr�{g�3UBRG���#ف]������m�<R���o!�[+S���AxP(u�l�%u��K���iŖP��=�ѫ׶E���J�r���fx����h���m�����` �B���H�OcGȕ���x29xRixG�u
�y<�~��U�o�m,��{i0 �HbCsg�g�O?���F!���!.N[~�˃�gQ�M�A�^wZET�jgp��"���6�2����(.42��
G�I�`�f����X˶l�����E���v҄n���`����[����q@ن�_MDS��/�T+�U�#���9&vv��
��t����?c���W�*��^?�m�˘��~�=ߟ�Y�V#�D�} =ۨ� �;i<3�/���ߒ������1����Yޗ���h�cqn[Z�A�#Pr-B?�'J9��b�����zXuj�_��5U=6U``-���'�b$ZJȄ��O���:#e���6���@`��G�s�Y���Ӎ��!�{�*L� �{�f�ͤo�E�n�R ]�׃�!0����2���K�Sꋑ�=�(V�T��P����/� ���r�%�x�JY��j��w��^!�S���SA�#U�W%�c3���
�h�-�fm�Zr��l@uW��q�Y�֖ݿ�5n��ǐ�;�i���JQ�2�+�OQ251r}B�Tލ�m�����;���XFD�d���NǝO ��r+W~d����Kn!P�i�rY��{]��p�h��M���Bz�Js(\�ZUX��rd(�繘z_P�o!�
=���[+w�z�W	�,����9�S��	�[%P�$@��h��R�{J���&^w����f��C/1,�~8]v���,�YS�re�0jx�;T�\;�J2���A���];���>߯AI�R珔�	LR�������(wu��@:���e��AT@0h��s'�RnK�܎��i�{���J�{~�9�A�>�x>Q���Ť�{�����聾����lW�4�t	"�R�
�A��(� �f �k	֛�d,��1�Ru���*�u����������|[7NڜvkE�~/'�t�V�c~����X�ɐ��?�~7w�j=/�&AU0�1�9^H��b�Y����^�R��{g�dWߚ�&���Ek���y���: 
��M�	N����~������F�Wex�`��6mó�xh��FK¼��m��z;�^/S[�x���B���?)2,e�~�uU�c�g�$)"?�����D�p�K��Njʄ	_��X���sC�G�Ds�� �^K���FEw&k�^��𻼁)����^s=���g�#|a������3?�6ˎ4j�\��m�+}*ԉX�D����U"�#l�虇;��vXx�K�f����i�w"���*֧��!w��/���L�k_p4�9)����nusfF��mV3������!������.o�ﵐ:\�  ��n~2{	M��澥'"q�*���<�����8�R��ܶ�0	�+ �V��ʨ��{ڏ����)�>?�b�F���w��O�?	E�n���6���վoo+�*)�]�JC_v�A6�����N������pQ>%��F��20V0E�w��;ǷJ74np* �1�;�?�?'�lC���Ψ���_<��A+�_���z#�n���I��������C��\��BP!�o]�}�黡ʜv7H�,�ip��禄tL�	�����h^�+U���t@�7*�Lā��BgL�iO��S�;Ɏ:��@^b[8�lQǑx��P�;�%nĔQ�-(�f���l���\�Q(���3�HЏy���!��'���o=��X8Y��_ٍ!�w:%�6�����3bGvf��:�,�r��=Z�q|X �7�N-�<:D��`�#	8�@bSG��)7�P�����\'du�^�ʌ]$�Gv9'����ݫG%��B�����Q�;�(�o�Ռ��8.I�����{�}���vcP\�ј��P��~�y���(n����Jǰ��oh�!��@��Z-3��ǯ_k('��叹��!Q�2j�/f���w�iz� �j`&{�������M� z6&�Q�����P �?dϬ@��PW`���w~B������ˢv\RZ�K����S%}Wo�A���
Q�[V�/�����|̯��K	ǵq�Gf���x��cޙTtǯ%N����ֺw�3��Ѩ2_�&�>Z��l���.eC�l�$W�^������b�Oȍ�����W�_)  K�_\\�����*C�jDb�Nr�y,�>j�O���+!g~�<F�'��)�>���`�A]>Б���k*�����Y�v��	��o]��>��@-�*�����{6U������N`��S��O�M�����=q#t��_�S�1�U�[�>X��l���%��r�����\�`���J�&p���K�'��R_�I�*b���Y�E�	��B���o�E։��:ݒF>D�py�`��M��6̳���6QH.��3�%o ������i�+��p|��� y
��\{�<���,t�Le*1�O�j�gz��	BBsŶqdj
8�	v��^o������U)�Cݖ����Һ����~��x�~
�d�h'�P!���R�\���˷��;��G�4#�����K�^�x�8����
�o�?s�yO{�r�`��Z�� J��d3�(�ƭ�
D�y��x��N�.��y�Dr���*.�Җ��.+T��Ϗ���N�_z�rB�����(���a3`��3�I��<PK0�ޒ:���K��0�M�Y%p?�����^��@�{��6��m8��?���Cړ`է�2�=y5�m�� k�R{�֐��=�������*A���dV����~N���HZ4�D&/�l#9����gt��:1���������O���3�OJKZ�'E��A]�[�� $��>�F4�Ls�7)������{.md�]�T(�w�x��:v���ѷzt�z+N�)I��!������E��C�H�P�}m�D��,7��+���>�\��uxٵFAX&F{��F����~��NR=��V��5����Z���UV8'v��,*c� vÛ�6W9�ofB�[_m�}2lK��4�6廹����=°ct�cC1B����m]{�a�\Z�Am���V�J,��Q ���.qJ���;�,�SN-�C��&��y��|к�3]픘����x�@Y�����%g�"��e&1����Jk�LbC��ԦD�b��V��|v�e��E3�0�y�a}��� �1ה͔gZ�Y�F�KԦ�呠�:��P��	��Dd�_�V��?2p��JR��`D5�{$���+�I��
@��ۘ�U��q�M�#z�X�k]$��¼���%Q5�1-�ol��Wg�jomd"ywI�dE�O�oPN�^�?6��ct���̇��ل�T?�Ӽw�L��/#��uI�m�D��dU�?��;���XL�,��Q�qa��̼�V����@N��6������1���GٙZ��y4&�iE�������dȦ����	��.a��y�BW�������>����i#W���#�_�,.��"�m7(D�"(�V�������d�t�1)&[S�Ҫ�����;�)Ɉ�)����ݡ:��t�[��jh�1�c��hɰ:�ϕl��b�:ȹ��$����j΍��A]�2&Q.C�.��2�FMnSg�����!�5T����&cT�Z�c���'y(�O���P����	�~���C��^��vj䄠g�	���h��vƥ�e<���;%Ɐ�Y��%V�k��!���L�g�����Ebb¨��e!퍓��uG$SS;�gU�� �4*���ʥ�
�? �bOC!�W��/Ł7@w���ػ�Tm����݈H�ƺ4:�nP��R*�m�@8s� W� r��u���o�JB2�쳉9���$��k���Pk��<N;"(�Ģ><�m���W�TŸߌ�yī0�َ��I�w<@���A4��`P5!���x��H㕧͆FwYF�}J>�]�)T�M ���@α��x(Å�g�=�����a�M�%���E^<�G��,p$H�,��Tz <l꘺������(��Q��;��Uql�M��.TZ�❀n�[h)�(w[���r���<yT\���K\��a�@�A�~%볗���h	߁^�*ɪ���j�m�MNN)!w�5%�X}��$B5[���0�1�4TT~��I-�%`�Չ�̛��c-ׇ�n��Iz�pr0Bf��3 �T�7A�3a�5A��M��6�iRN��o�}�f���k���.cu|�F#ؾp�Z���,-�!����O t��t���j���k�^XB5���>��F������>>[�o����OL�Ȫ�?�F��@�ܜ�<0�7�@~�-3A�c ��m�ge����0i��BZ��A9�BW