��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�M�N��.��	F(�
F[)b��5!�J��}F���Iu#:z�ϫD[H�LnΦ��w!��j�k�tBB(&b.��Y��,b�)�{������Z��-�C̷/��0Hm��a�
� �?�#�^�Oim1�3��b�qÁ�@9d�5���|H{�S�/!�K���z�<��d�,�I��C�3�B0�%��mKv�nJ��Z	WT\ЇHڲ.�ѻx�w���/�u+]�b��X(TVŇ��L���a�6{����bka�$z4����ߟ;Q?�^���v��I����y�~�#��-P�d$��a��H�$P?�R������-�b?*���Ɓq��.v�
C��8�t�m���q>�K�(f<&�o{8�������4��9&WǗT��Ƨ9����Þ�����ò�$�(ʘ�4݇�Y�	���#&Ce=4؉(����� �w�{C>;7�L��)Ĭ*$���ձA!����I��/
#�{>�"zm]7���w���Ͻ��%��6�y�=�i	x�jQgW�N�}~���cS��Ne���4�
Ӡ$
K�D
���t]2)e�+_����f&�@��h�U��h<����X��*��{��z8�$�b�\̑��.���A���:=���ɯ�lu��2[��1�l�?qW7�?(����:p] ����v��Ng]7^��.&��i�x�z��� J��\) ��;�a�Y8u�G�l��w�%��r��ݟ0
BW�����@�[+�:�:Ǿ��Z©�WQh��Ϥ�`�.~3��ɣ^�ґn�*#��Z��;g�|+F5+I���\�Ǝ���0ĵ��/G.���JS\
0Zw3�L��`�M��`q!�Ís�L��֕���(7*sG�V$�=�{T����qc�B��ޮ����F�k10����V��7��i�/H�G%��Z>�adZ%����м:Y�2��u���4Zۇ1��_=f$q��y����g0N��;�#�P˄_�o75�G�೷�0����+�&��8���P�L�Z3���C/}��Q0u������>7Չt��J����?����r�]���w*)��=����s���ŚT�=��bѬ5�A�R�Q\d��t�5e$�v��h �IG-����R~�cR4;���H�]��I-BF��p+����8� ���
Z��5���� �ܦ��s=icw�$�3?�{��W��V���2��:" 睷LA��I���t��*$N�f�p��g�f��&L���P���~r���-���A�TEl���1ǩ������׉T�u/���u��8mI�w.Z�Yf����"Z�Ŋ��xр�\����i�6QtP}��Яˁ�*��r��<�/Y��g��(Q�O7݉��RV�y�(R^|vÂg�'��G���F%��ª������Zۓlx;���P�ʫ�L��0V5��X��� �|��ˈ�NN%��	$�B��!���W��S���D��M�]�b�	?�du��\\�a2��`�n�Vt�l��nE�7�vw&^<���	j��ҭe��P�誄�*�(��G��4�M*D�
� pY�ڳ���rd�T���yv��.E�*s�/Sl5E�'Tt�`�_�}&0)mXt��0���ݦ9�E[_:.@z/S��Ɗ4u���H+��a���ݱ`���]ۯ���m�8-�e$��X���HkJ�#�d�Gg!V�a3�F����(�I[��=V�)<��El%Վ�G|/�-����A��*?���l �^���7��D2�y�:�;C�p ��?Hݤi�㰐gӘ���ڿ4���툭��� �x�M^W>�tt��=�Z���	�Lr*������,:|0|d<S�Y�0�4��~��v��9��;��S���Va�'@W�b!�Nο��\N��k*�䉗!:"T�f���A�=�1D�:�!7S�J��11^\�����^}��)��ʴ�pu��7��������U�����9<����Q�OZ�d>�Hib�0�b;���3(������	:�*�.�Z�;{�1���h���a�AtOO��.0�ȓa������7�K��Ϸ�x�,}�K��;��58�Z�$U�xz��l�J+4�ꋌ#zO�I5�6̠���ސO'g$�g�Pw�i
�4�lXri����N)����.-�UA�4�o����[���uĬ�<]p����%���:�z&U�{�sޒ�Mɳ8i�W:(�_Իn)`�M�Ʊr/����r�d��N�	ל��^;)���D�+�C��[�#�@�>זx�
��Z�G'Ԫ�=C�@ۜ2�c�s��(	D
�-G�i�|q|4P�D4���"�s��rr�N�w�ML�Q?�Gh$�����}G���P��ʒk54@F�g����M��?Ձ#'�ȅ��r�Y��$�g�u�o�Ee�����FP�6�ԳEc�������3��3�%�L��{�x���*�2�+�P&@v?f����������E��i�;��#<�1��f_�%dM�_��V�RV;��F��-'�dg6Aŋ,n�T<Z�֓�?��+KY��ynx�����_XQx�J�-�Ӯ{E<}7��^EvV�%mbݨ�����(����j�L ���(�Ԑ}�	�d�foD �����(���wള�X�d���~n���«=i�M�F���Vi��-��l_�5b�](��,@��1��;
��cyK��s�5g��7�
�w�d�����������ԨMq����N�՝�Q�s<z����M�n��0}���~�M�,���B���q�}l���ӱ:S����0?��DW�X�@>��q��Fl3a��w�������V,G���ʹKq���?�0��8-��N5�g@Ŝ/+k�M'*�i��qP����X�/�#��w��((�8�SkӈI�(�sd<�k����=Ͽ���&�A;/��Y$N��;TL�oj@q�9w���*�!�>�i���i���X��cB�ٓ�(�;P�p�I�(�G�5��oe������g�\�@��J�`�z��ύ��8�}�	7fȕɴ���w>�����;p^�iin�w�N����8�gqP���C�5��
gB0�y���p�̀�"����U&_��e8��f_`�1Wy��ڹ�Ie���z�e��ʑ�N�A&��}�8BӾ.�r[�t:�qm<�_��"��>a���2!�	lT�^���z��mOB��~
f�-���y�B��y�e����-�CAĶKht��-l&��`�w�r&�h���b�Ng;km�$ވJ(����G*%?�K�߁��b��ެH���i����v�֙0,k~u�l��c����پ9gJ;?�E��䦤�Ƞ�|���q\��S��4gtڋ!:W4\��ٗ�x��B���\���M�s���awu�/��Ԗ�]����ҙan�F�����q��Yg�n��PHk$���t�2qp=N�@�g{=��O�*�b�4��V&��1�~~:nk����ky��1�v�h$O�t����._>C�+i���,�V)Jć�FFVx�Q���_#Y�9�Jd>�S%�� I��\�?y���Ȑ4χ8ٺ���x��J�Xc��%�}W�r� �9?X��TC�� rQ��D~R3�\�KBH+�q�O��#z�y.ߕx����!?��v�'[�[�/��;?���b	ybX
��{wI�켎?���QU-=i
˿�ׂ�*_�+��쒏g
�j�YЙ����5n����tr���8�g�JA`(E��P��+�AM�6�NP-n��"qq+��둮�=�"�hZ�7�.�(�z���z��G߻	�9M���\LB��9�Zh�)p V�]J=>Ƌ8	&`2�zo�����[���%*�."�,��2Oz�_��t�N�U' ��9ң�<��U�'у�4�ɒV��qJ�����e���1������CH"��zq�8��[#�ˀ�P��y���^/�k��R�-ئAje�Ή�u�o7�:E��կ�4���oB��f��PS3}�v�Y��֕_�����tIL5y�u��>��W���ϧ��H�l?�"����L�t��p���2�b]�y<Ĵ5)jx��$�x��1�
D_͜�P�?C����~�p�o����#�m�Ҡ����|	]�a��<3e��>�,�ZPM�<7�"ɐ�I��#��J�O���)�e�"���@m��HqS��?�NRSt"����lh֨9eG�